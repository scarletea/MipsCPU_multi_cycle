module EXT(
   input  [15:0] Imm16,
   input  [1:0]  EXTOp,
   output reg [31:0] Imm32
};
